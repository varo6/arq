library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity programa_helloworld_int_FLIP is
	port( address : in std_logic_vector(15 downto 0);
		clk : in std_logic;
		dout : out std_logic_vector(25 downto 0));
	end;

architecture v1 of programa_helloworld_int_FLIP is

	constant ROM_WIDTH: INTEGER:= 26;
	constant ROM_LENGTH: INTEGER:= 65536;

	subtype rom_word is std_logic_vector(ROM_WIDTH-1 downto 0);
	type rom_table is array (0 to ROM_LENGTH-1) of rom_word;

constant rom: rom_table := rom_table'(
	"01111000000000000000000000",
	"01101100000000000000001111",
	"00000001110000000000000000",
	"01100011000111000000000000",
	"00010011000000000000000000",
	"01101010000000000000001001",
	"01101100000000000000011100",
	"00010001110000000000000001",
	"01101000000000000000000011",
	"01111000000000000000000001",
	"00000001100000000000001001",
	"00011001100000000000000001",
	"01101010100000000000001011",
	"00000001100000000000001001",
	"01101000000000000000001011",
	"01000010000000000011111111",
	"00000110001000000000000000",
	"01101010100000000000001111",
	"01101100000000000000110000",
	"00000000110000000000010001",
	"01101100000000000000101001",
	"01010010000000000000001110",
	"01000000000000000011111111",
	"00000100001000000000000000",
	"00101010000000000000000000",
	"00011000110000000000000001",
	"01101010100000000000010100",
	"01001000000000000000000000",
	"00000000000000000000000000",
	"01000100000000000011111111",
	"01101100000000000000101001",
	"00000000110000000000001000",
	"01000111000000000011111111",
	"01101100000000000000101001",
	"01010011000000000000001110",
	"00011000110000000000000001",
	"01101010100000000000100000",
	"00000000000000000011111111",
	"01000100000000000011111111",
	"01101100000000000000101001",
	"01001000000000000000000000",
	"00000001000000000000000011",
	"00000001010000000000100010",
	"00011001010000000000000001",
	"01101010100000000000101011",
	"00011001000000000000000001",
	"01101010100000000000101010",
	"01001000000000000000000000",
	"00000001000000000000000011",
	"00000001010000000000010000",
	"00011001010000000000000001",
	"01101010100000000000110010",
	"00011001000000000000000001",
	"01101010100000000000110001",
	"01001000000000000000000000",
	"01111000000000000000000000",
	"01101100000000000000001111",
	"00100011001000000000000000",
	"01101100000000000000011100",
	"00010001100000000000110000",
	"00100011000110000000000000",
	"01101100000000000000011100",
	"01011000000000000000000001",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"01101000000000000000110111");

begin

process (clk)
begin
	if clk'event and clk = '1' then
		dout <= rom(conv_integer(address));
	end if;
end process;
end v1;
