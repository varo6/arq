library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity programa_helloworld_int_FLIP is
	port( address : in std_logic_vector(7 downto 0);
		clk : in std_logic;
		dout : out std_logic_vector(15 downto 0));
	end;

architecture v1 of programa_helloworld_int_FLIP is

	constant ROM_WIDTH: INTEGER:= 16;
	constant ROM_LENGTH: INTEGER:= 256;

	subtype rom_word is std_logic_vector(ROM_WIDTH-1 downto 0);
	type rom_table is array (0 to ROM_LENGTH-1) of rom_word;

constant rom: rom_table := rom_table'(
	"1111000000000000",
	"1101100000001111",
	"0000011100000000",
	"1100000111100000",
	"0010000100000000",
	"1101010000001001",
	"1101100000011100",
	"0010011100000001",
	"1101000000000011",
	"1111000000000001",
	"0000011000001001",
	"0011011000000001",
	"1101010100001011",
	"0000011000001001",
	"1101000000001011",
	"1000001011111111",
	"0000101010000000",
	"1101010100001111",
	"1101100000110000",
	"0000001100001001",
	"1101100000101001",
	"1010001000001110",
	"1000000011111111",
	"0000100010000000",
	"0101001000000000",
	"0011001100000001",
	"1101010100010100",
	"1001000000000000",
	"0000000000000000",
	"1000100011111111",
	"1101100000101001",
	"0000001100001000",
	"1000100111111111",
	"1101100000101001",
	"1010000100001110",
	"0011001100000001",
	"1101010100100000",
	"0000000011111111",
	"1000100011111111",
	"1101100000101001",
	"1001000000000000",
	"0000010000000011",
	"0000010100100010",
	"0011010100000001",
	"1101010100101011",
	"0011010000000001",
	"1101010100101010",
	"1001000000000000",
	"0000010000000011",
	"0000010100010000",
	"0011010100000001",
	"1101010100110010",
	"0011010000000001",
	"1101010100110001",
	"1001000000000000",
	"1111000000000000",
	"1101100000001111",
	"1111101000000000",
	"0100000101000000",
	"1101100000011100",
	"0010011000110000",
	"0100000111000000",
	"1101100000011100",
	"1011000000000001",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"1101000000110111");

begin

process (clk)
begin
	if clk'event and clk = '1' then
		dout <= rom(conv_integer(address));
	end if;
end process;
end v1;
