library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity test_instrucciones is
	port( address : in std_logic_vector(15 downto 0);
		clk : in std_logic;
		dout : out std_logic_vector(25 downto 0));
	end;

architecture v1 of test_instrucciones is

	constant ROM_WIDTH: INTEGER:= 26;
	constant ROM_LENGTH: INTEGER:= 65536;

	subtype rom_word is std_logic_vector(ROM_WIDTH-1 downto 0);
	type rom_table is array (0 to ROM_LENGTH-1) of rom_word;

constant rom: rom_table := rom_table'(
	"11010000000000000000001111",
	"11010010000000000000001111",
	"11010010100000000000001111",
	"11010011000000000000001111",
	"11010011100000000000001111",
	"11011000000000000000001111",
	"11011010000000000000001111",
	"11011010100000000000001111",
	"11011011000000000000001111",
	"11011011100000000000001111",
	"10010000000000000000000000",
	"10010010000000000000000000",
	"10010010100000000000000000",
	"10010011000000000000000000",
	"10010011100000000000000000",
	"10100011110000000000001110",
	"10100010010000000000001111",
	"10100010010000000000001010",
	"10100010010000000000001000",
	"10100010010000000000001100",
	"10100010010000000000000110",
	"10100010010000000000000111",
	"10100010010000000000000010",
	"10100010010000000000000000",
	"10100010010000000000000100",
	"00000010101011011111100000",
	"00001010101011011111100000",
	"00010010101011011111100000",
	"00011010101011011111100000",
	"01000010101111000000000000",
	"01001010101111000000000000",
	"01010010101111000000000000",
	"01011010101111000000000000",
	"00100011101011011111100000",
	"00101011101011011111100000",
	"00110011101011011111100000",
	"00111011101011011111100000",
	"01100011101011000000000000",
	"01101011101011000000000000",
	"01110011101011000000000000",
	"01111011101011000000000000",
	"10000010001011010110010111",
	"11000010001100000000000000",
	"10001010001011010110010111",
	"11001010001100000000000000",
	"11110000000000000000000001",
	"11110000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000",
	"00000000000000000000000000");

begin

process (clk)
begin
	if clk'event and clk = '1' then
		dout <= rom(conv_integer(address));
	end if;
end process;
end v1;
