library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity programa_ahorcado is
	port( address : in std_logic_vector(7 downto 0);
		clk : in std_logic;
		dout : out std_logic_vector(15 downto 0));
	end;

architecture v1 of programa_ahorcado is

	constant ROM_WIDTH: INTEGER:= 16;
	constant ROM_LENGTH: INTEGER:= 256;

	subtype rom_word is std_logic_vector(ROM_WIDTH-1 downto 0);
	type rom_table is array (0 to ROM_LENGTH-1) of rom_word;

constant rom: rom_table := rom_table'(
	"1111000000000000",
	"1101100000000100",
	"1111000000000001",
	"1101000000000001",
	"1000001011111111",
	"0000101010000000",
	"1101010100000100",
	"1101100000100101",
	"0000001100001001",
	"1101100000011110",
	"1010001000001110",
	"1000000011111111",
	"0000100010000000",
	"0101001000000000",
	"0011001100000001",
	"1101010100001001",
	"1001000000000000",
	"0000000000000000",
	"1000100011111111",
	"1101100000011110",
	"0000001100001000",
	"1000100111111111",
	"1101100000011110",
	"1010000100001110",
	"0011001100000001",
	"1101010100010101",
	"0000000011111111",
	"1000100011111111",
	"1101100000011110",
	"1001000000000000",
	"0000010000000011",
	"0000010100100010",
	"0011010100000001",
	"1101010100100000",
	"0011010000000001",
	"1101010100011111",
	"1001000000000000",
	"0000010000000011",
	"0000010100010000",
	"0011010100000001",
	"1101010100100111",
	"0011010000000001",
	"1101010100100110",
	"1001000000000000",
	"0000011000000000",
	"1100000111000000",
	"0010000100000000",
	"1101010000110011",
	"1101100000010001",
	"0010011000000001",
	"1101000000101101",
	"1001000000000000",
	"0000000100001010",
	"1101100000010001",
	"0000000100001101",
	"1101100000010001",
	"0000000101001100",
	"1101100000010001",
	"0000000101000101",
	"1101100000010001",
	"0000000101010100",
	"1101100000010001",
	"0000000101010010",
	"1101100000010001",
	"0000000101000001",
	"1101100000010001",
	"0000000100111010",
	"1101100000010001",
	"0000000100100000",
	"1101100000010001",
	"1001000000000000",
	"0000000100001010",
	"1101100000010001",
	"0000000100001101",
	"1101100000010001",
	"0000000101010010",
	"1101100000010001",
	"0000000101000101",
	"1101100000010001",
	"0000000100111010",
	"1101100000010001",
	"0000000100100000",
	"1101100000010001",
	"1001000000000000",
	"0000000100001010",
	"1101100000010001",
	"0000000100001101",
	"1101100000010001",
	"0000000101001101",
	"1101100000010001",
	"0000000101010101",
	"1101100000010001",
	"0000000101000011",
	"1101100000010001",
	"0000000101001000",
	"1101100000010001",
	"0000000101001111",
	"1101100000010001",
	"0000000101010011",
	"1101100000010001",
	"0000000100100000",
	"1101100000010001",
	"0000000101000101",
	"1101100000010001",
	"0000000101010010",
	"1101100000010001",
	"0000000101010010",
	"1101100000010001",
	"0000000101001111",
	"1101100000010001",
	"0000000101010010",
	"1101100000010001",
	"0000000101000101",
	"1101100000010001",
	"0000000101010011",
	"1101100000010001",
	"0000000100100001",
	"1101100000010001",
	"1101000000000001",
	"0000000100001010",
	"1101100000010001",
	"0000000100001101",
	"1101100000010001",
	"0000000101010111",
	"1101100000010001",
	"0000000101001001",
	"1101100000010001",
	"0000000101001110",
	"1101100000010001",
	"0000000100100001",
	"1101100000010001",
	"1101000000000001",
	"0000000100001010",
	"1101100000010001",
	"0000000100001101",
	"1101100000010001",
	"0000000101000101",
	"1101100000010001",
	"0000000101010010",
	"1101100000010001",
	"0000000101010010",
	"1101100000010001",
	"0000000101001111",
	"1101100000010001",
	"0000000101010010",
	"1101100000010001",
	"0000000101000101",
	"1101100000010001",
	"0000000101010011",
	"1101100000010001",
	"0000000100111010",
	"1101100000010001",
	"0000000100100000",
	"1101100000010001",
	"1000011101001001",
	"0100000111100000",
	"0010000100110000",
	"1101100000010001",
	"1001000000000000",
	"1000011101001001",
	"1101100010000100",
	"0100011011100000",
	"0011011000001001",
	"1101011101010100",
	"1101000010100101",
	"1101100000110100",
	"1101100000000100",
	"0100000101000000",
	"1101100000010001",
	"1000101001000101",
	"1101100000011110",
	"1000101001000110",
	"1101100001000111",
	"1000000101000110",
	"1000100101000111",
	"1111100100000000",
	"0100011000100000",
	"1101100000010001",
	"0001111001000110",
	"1101010001110111",
	"1101000010011111",
	"1111000000000000",
	"0000000100000000",
	"1101100000101100",
	"1101100000011110",
	"1101100000011110",
	"1101100000000100",
	"1000101001000001",
	"1101100000011110",
	"1101100000000100",
	"1000101001000010",
	"1101100000011110",
	"1101100000000100",
	"1000101001000011",
	"1101100000011110",
	"1101100000000100",
	"1000101001000100",
	"1101100000011110",
	"1101000010100101",
	"1011000000000001",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"0000000000000000",
	"1101000010110101");

begin

process (clk)
begin
	if clk'event and clk = '1' then
		dout <= rom(conv_integer(address));
	end if;
end process;
end v1;
